module controller #(parameter SIZE = 32) (
	input clk,
	output read,
	output reg en_S2, en_C3, en_S4, en_C5
);

endmodule
